/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */
`default_nettype none
`timescale 1ns / 1ps

module tt_um_fifo #(parameter DSIZE=8, parameter ASIZE=4) (
    input  wire [7:0]  ui_in,    // Switches (input data)
    output wire [7:0]  uo_out,   // LEDs (read data output)
    input  wire [7:0]  uio_in,   // IOs: Input path (write/read control & resets)
    output wire [7:0]  uio_out,  // IOs: Output status path (flags, clocks)
    output wire [7:0]  uio_oe,   // IOs: Output enable path (active high: output, else input)
    input  wire        ena,      // Enable (always 1 on Tiny Tapeout platform)
    input  wire        clk,      // 100 MHz system clock
    input  wire        rst_n     // Global reset (active low)
);

    // Assign write/read control and reset from IO inputs
    wire winc = uio_in[7];      // Write increment enable
    wire rinc = uio_in[6];      // Read increment enable
    wire rrst_n = uio_in[3];    // Read side reset (active low)
    wire wrst_n = uio_in[4];    // Write side reset (active low)

    // Write and read data buses
    wire [DSIZE-1:0] wdata = ui_in;
    wire [DSIZE-1:0] rdata;

    // Full and empty signals
    wire wfull, rempty;

    // Internal clocks generated by clock divider
    wire wclk, rclk;

    // Assign always-on output enable signals for the IO output pins where needed
    // Output enables: 1=drive output, 0=high-z/input mode
    assign uio_oe = 8'b00100111; // Bits 0,1,2,4,5 driven as output

    // Drive status flags and clocks onto IO output pins
    assign uio_out[0] = rempty;  // FIFO empty status
    assign uio_out[1] = wfull;   // FIFO full status
    assign uio_out[2] = rclk;    // Read clock
    assign uio_out[5] = wclk;    // Write clock

    // Drive zeros to unused output bits
    assign uio_out[7:6] = 2'b00;
    assign uio_out[4:3] = 2'b00;

    // Output read data to LEDs
    assign uo_out = rdata;

    // Clock divider instance to create asynchronous clocks
    clock_div clk_div_inst (
        .clk   (clk),
        .rst_n (rst_n),
        .wclk  (wclk),
        .rclk  (rclk)
    );

    // Pointer synchronization wires
    wire [ASIZE:0] wptr, rptr;
    wire [ASIZE:0] WSR2_ptr, RSW2_ptr;

    // Write enable and read enable signals gated with full and empty flags
    wire wclken = (winc && !wfull);
    wire rclken = (rinc && !rempty);

    // Synchronizers for crossing clock domains - read to write pointer sync
    sync_R2W sync_r2w (
        .RSW2_ptr(RSW2_ptr),
        .rptr(rptr),
        .wclk(wclk),
        .wrst_n(wrst_n)
    );

    // Synchronizers for crossing clock domains - write to read pointer sync
    sync_W2R sync_w2r (
        .WSR2_ptr(WSR2_ptr),
        .wptr(wptr),
        .rclk(rclk),
        .rrst_n(rrst_n)
    );

    // FIFO memory block instance
    fifomem #(DSIZE, ASIZE) fifomem_inst (
        .rdata(rdata),
        .wdata(wdata),
        .raddr(rptr[ASIZE-1:0]),
        .waddr(wptr[ASIZE-1:0]),
        .wclken(wclken),
        .wclk(wclk),
        .rclken(rclken),
        .rclk(rclk)
    );

    // Empty flag and read pointer management
    rptr_empty #(.ASIZE(ASIZE)) rptr_empty_inst (
        .rempty(rempty),
        .raddr(rptr[ASIZE-1:0]),
        .rptr(rptr),
        .WSR2_ptr(WSR2_ptr),
        .rinc(rinc),
        .rclk(rclk),
        .rrst_n(rrst_n)
    );

    // Full flag and write pointer management
    wptr_full #(.ASIZE(ASIZE)) wptr_full_inst (
        .wfull(wfull),
        .waddr(wptr[ASIZE-1:0]),
        .wptr(wptr),
        .RSW2_ptr(RSW2_ptr),
        .winc(winc),
        .wclk(wclk),
        .wrst_n(wrst_n)
    );

    // Use all unused inputs to prevent synthesis warnings
    wire _unused = &{ena, uio_in[5], uio_in[2:0], rst_n};

endmodule
